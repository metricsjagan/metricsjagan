package ahb_master_agent_pkg;

import uvm_pkg::*;
  //`include "uvm_macros.svh"



  `include "ahb_master_defines.sv"
  `include "ahb_master_types.sv"
  `include "ahb_master_transaction_c.sv"

  `include "ahb_master_sequencer.sv"
  `include "ahb_master_driver.sv"
  `include "ahb_master_monitor.sv"
  `include "ahb_master_agent_config.sv"
  `include "ahb_master_agent.sv"


endpackage: ahb_mater_agent_pkg
