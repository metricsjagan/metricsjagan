module tb_top();
  
  input [31:0] haddr;
  input        hmastlock;
  input [2:0]  hsize;
  input [1:0]  htrans;
  input [31:0] hwdata;
  input        hwrite;
  output [31:0] hrata;
  output        hready;
  output       hresp;
  
  
  
  
  
  
  
endmodule 
